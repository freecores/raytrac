--! @file raytrac.vhd
--! @brief Descripci�n del sistema aritmetico usado por raytrac.
--! @author Juli�n Andr�s Guar�n Reyes.
-- RAYTRAC
-- Author Julian Andres Guarin
-- uf.vhd
-- This file is part of raytrac.
-- 
--     raytrac is free software: you can redistribute it and/or modify
--     it under the terms of the GNU General Public License as published by
--     the Free Software Foundation, either version 3 of the License, or
--     (at your option) any later version.
-- 
--     raytrac is distributed in the hope that it will be useful,
--     but WITHOUT ANY WARRANTY; without even the implied warranty of
--     MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
--     GNU General Public License for more details.
-- 
--     You should have received a copy of the GNU General Public License
--     along with raytrac.  If not, see <http://www.gnu.org/licenses/>.

--! Libreria de definicion de senales y tipos estandares, comportamiento de operadores aritmeticos y logicos.\n Signal and types definition library. This library also defines 
library ieee;
--! Paquete de definicion estandard de logica. Standard logic definition pack.
use ieee.std_logic_1164.all;
--! Se usaran en esta descripcion los componentes del package arithpack.vhd.\n It will be used in this description the components on the arithpack.vhd package. 
use work.arithpack.all;


--! uf es la descripci�n del circuito que realiza la aritm�tica del Rt Engine.

--! La entrada opcode indica la operaci�n que se est� realizando, en los sumadores, es la misma se�al que se encuentra en la entidad opcoder, que selecciona si se est� realizando un producto punto o un producto cruz. Dentro de la arquitectura de uf, la se�al opcode selecciona en la primera etapa de sumadores, si la operaci�n a realizar ser� una resta o una suma. 
--! Los resultados estar�n en distintas salidas dependiendo de la operaci�n, lo cual es apenas natural: El producto cruz tiene por resultado un vector, mientras que el producto punto tiene por resultado un escalar. 
--! Esta entidad utiliza las se�ales de control clk y rst.}
--! \n\n
--! La caracter�stica fundamental de uf, es que puede realizar 2 operaciones de producto punto al mimso tiempo � una operaci�n de producto cruz al mismo tiempo. La otra caracter�stica importante es que el pipe de producto punto es mas largo que el pipe de producto cruz: el producto punto tomar� 3 clocks para realizarse, mientras que el procto punto tomara 4 clocks para realizarse.    

entity uf is 
	port (
		opcode		: in std_logic; --! Entrada que dentro de la arquitectura funciona como selector de la operaci�n que se lleva a cabo en la primera etapa de sumadores/restadores. 
		m0f0,m0f1,m1f0,m1f1,m2f0,m2f1,m3f0,m3f1,m4f0,m4f1,m5f0,m5f1 : in std_logic_vector(17 downto 0); --! Entradas que van conectadas a los multiplicadores en la primera etapa de la descripci�n.  
		cpx,cpy,cpz,dp0,dp1 : out std_logic_vector(31 downto 0); --! Salidas donde se registran los resultados de las operaciones aritm�ticas: cpx,cpy,cpz ser�n los componentes del vector que da por resultado el producto cruz entre los vectores AxB � CxD.  
		clk,rst		: in std_logic --! Las entradas de control usuales.  
	);
end uf;

architecture uf_arch of uf is 

	-- Stage 0 signals
	
	signal stage0mf00,stage0mf01,stage0mf10,stage0mf11,stage0mf20,stage0mf21,stage0mf30,stage0mf31,stage0mf40,stage0mf41,stage0mf50,stage0mf51 : std_logic_vector(17 downto 0); --! Se�ales que conectan los operandos seleccionados en opcode a las entradas de los multiplicadores.
	signal stage0p0,stage0p1, stage0p2, stage0p3, stage0p4, stage0p5 : std_logic_vector(31 downto 0); --! Se�ales / buses, con los productos de los multiplicadores. 
	signal stage0opcode : std_logic; --! Se�al de atraso del opcode. Revisar el diagrama de bloques para mayor claridad.
	
	--Stage 1 signals 
	
	signal stage1p0, stage1p1, stage1p2, stage1p3, stage1p4, stage1p5 : std_logic_vector (31 downto 0); --! Se�ales provenientes de los productos de la etapa previa de multiplicadores.
	signal stage1a0, stage1a1, stage1a2 : std_logic_vector (31 downto 0); --! Se�ales / buses, con los resultados de los sumadores. 
	signal stage1opcode : std_logic; --! Se�al proveniente del opcode que selecciona si los sumadores deben ejecutar una resta o una suma dependiendo de la operaci�n que se ejecute en ese momento del pipe.  
	
	-- Some support signals
	signal stage1_internalCarry	: std_logic_vector(2 downto 0); --! Cada uno de los 3 sumadores de la etapa de sumadores est� compuesto de una cascada de 2 sumadores Carry Look Ahead: aXhigh y aXlow. El carry out del componente low y el carry in del componente high, se conectar� a trav�s de las se�ales internal carry.   
	signal stage2_internalCarry : std_logic_vector(1 downto 0); --! Cada uno de los 2 sumadores de la �ltima etapa de sumadores est� compuesto de una cascada de 2 sumadores Carry Look Ahead�: aXhigh y aXlow. El carry out del componente low y el carry in del componente high, se conectar� a trav�s de las se�ales internal carry.  
	
	--Stage 2 signals	
	signal stage2a0, stage2a2, stage2a3, stage2a4, stage2p2, stage2p3 : std_logic_vector (31 downto 0); --! Estas se�ales corresponden a los sumandos derivados de la primera etapa de multiplicadores (stage2p2, stage2p3) y a los sumandos derivados del resultado de las sumas en la primera etapa de sumadores. 
	
	  	
	
begin

	-- Multiplicator Instantiation (StAgE 0)
	--! Multiplicador 0 
	m0 : r_a18_b18_smul_c32_r 
	port map (
		aclr	=> rst,
		clock	=> clk,
		dataa	=> stage0mf00,
		datab	=> stage0mf01,
		result	=> stage0p0
	);
	
	--! Multiplicador 1
	m1 : r_a18_b18_smul_c32_r 
	port map (
		aclr	=> rst,
		clock	=> clk,
		dataa	=> stage0mf10,
		datab	=> stage0mf11,
		result	=> stage0p1
	);
	
	--! Multiplicador 2
	m2 : r_a18_b18_smul_c32_r 
	port map (
		aclr	=> rst,
		clock	=> clk,
		dataa	=> stage0mf20,
		datab	=> stage0mf21,
		result	=> stage0p2
	);
	
	--! Multiplicador 3
	m3 : r_a18_b18_smul_c32_r 
	port map (
		aclr	=> rst,
		clock	=> clk,
		dataa	=> stage0mf30,
		datab	=> stage0mf31,
		result	=> stage0p3
	);
	
	--! Multiplicador 4
	m4 : r_a18_b18_smul_c32_r 
	port map (
		aclr	=> rst,
		clock	=> clk,
		dataa	=> stage0mf40,
		datab	=> stage0mf41,
		result	=> stage0p4
	);
	
	--! Multiplicador 5
	m5 : r_a18_b18_smul_c32_r 
	port map (
		aclr	=> rst,
		clock	=> clk,
		dataa	=> stage0mf50,
		datab	=> stage0mf51,
		result	=> stage0p5
	);
	
	-- Adder Instantiation (sTaGe 1)
	
	--! Adder 0, 16 bit carry lookahead low adder. 
	a0low : adder 
	generic map (
		16,"CLA","YES"	-- Carry Look Ahead Logic (More Gates Used, But Less Time)
						-- Yes instantiate Xor gates stage in the adder so we can substract on the opcode signal command.
	)
	port map	(
		a => stage1p0(15 downto 0),
		b => stage1p1(15 downto 0),
		s => stage1opcode,
		ci => '0',
		result => stage1a0(15 downto 0),
		cout =>	stage1_internalCarry(0)
	);
	--Adder 0, 16 bit carry lookahead high adder.
	a0high : adder 
	generic map (
		w => 16,
		carry_logic 		=> "CLA",	-- Carry Look Ahead Logic (More Gates Used, But Less Time)
		substractor_selector	=> "YES"	-- Yes instantiate Xor gates stage in the adder so we can substract on the opcode signal command.
	)
	port map	(
		a => stage1p0(31 downto 16),
		b => stage1p1(31 downto 16),
		s => stage1opcode,
		ci => stage1_internalCarry(0),
		result => stage1a0(31 downto 16),
		cout =>	open
	);
	--! Adder 1, 16 bit carry lookahead low adder. 
	a1low : adder 
	generic map (
		w => 16,
		carry_logic 		=> "CLA",	-- Carry Look Ahead Logic (More Gates Used, But Less Time)
		substractor_selector	=> "YES"	-- Yes instantiate Xor gates stage in the adder so we can substract on the opcode signal command.
	)
	port map	(
		a => stage1p2(15 downto 0),
		b => stage1p3(15 downto 0),
		s => stage1opcode,
		ci => '0',
		result => stage1a1(15 downto 0),
		cout =>	stage1_internalCarry(1)
	);
	--! Adder 1, 16 bit carry lookahead high adder.
	a1high : adder 
	generic map (
		w => 16,
		carry_logic 		=> "CLA",	-- Carry Look Ahead Logic (More Gates Used, But Less Time)
		substractor_selector	=> "YES"	-- Yes instantiate Xor gates stage in the adder so we can substract on the opcode signal command.
	)
	port map	(
		a => stage1p2(31 downto 16),
		b => stage1p3(31 downto 16),
		s => stage1opcode,
		ci => stage1_internalCarry(1),
		result => stage1a1(31 downto 16),
		cout =>	open
	);	
	--! Adder 2, 16 bit carry lookahead low adder. 
	a2low : adder 
	generic map (
		w => 16,
		carry_logic 		=> "CLA",	-- Carry Look Ahead Logic (More Gates Used, But Less Time)
		substractor_selector	=> "YES"	-- Yes instantiate Xor gates stage in the adder so we can substract on the opcode signal command.
	)
	port map	(
		a => stage1p4(15 downto 0),
		b => stage1p5(15 downto 0),
		s => stage1opcode,
		ci => '0',
		result => stage1a2(15 downto 0),
		cout =>	stage1_internalCarry(2)
	);
	--! Adder 2, 16 bit carry lookahead high adder.
	a2high : adder 
	generic map (
		w => 16,
		carry_logic 		=> "CLA",	-- Carry Look Ahead Logic (More Gates Used, But Less Time)
		substractor_selector	=> "YES"	-- Yes instantiate Xor gates stage in the adder so we can substract on the opcode signal command.
	)
	port map	(
		a => stage1p4(31 downto 16),
		b => stage1p5(31 downto 16),
		s => stage1opcode,
		ci => stage1_internalCarry(2),
		result => stage1a2(31 downto 16),
		cout =>	open
	);
	
	
	-- Adder Instantiation (Stage 2)
	--! Adder 3, 16 bit carry lookahead low adder. 
	a3low : adder 
	generic map (
		w => 16,
		carry_logic 		=> "CLA",	-- Carry Look Ahead Logic (More Gates Used, But Less Time)
		substractor_selector	=> "NO"		-- No Just Add.
	)
	port map	(
		a => stage2a0(15 downto 0),
		b => stage2p2(15 downto 0),
		s => '0',
		ci => '0',
		result => stage2a3(15 downto 0),
		cout =>	stage2_internalCarry(0)
	);
	--Adder 3, 16 bit carry lookahead high adder.
	a3high : adder 
	generic map (
		w => 16,
		carry_logic 		=> "CLA",	-- Carry Look Ahead Logic (More Gates Used, But Less Time)
		substractor_selector	=> "NO"		-- No Just Add.
	)
	port map	(
		a => stage2a0(31 downto 16),
		b => stage2p2(31 downto 16),
		s => '0',
		ci => stage2_internalCarry(0),
		result => stage2a3(31 downto 16),
		cout =>	open
	);
	--! Adder 4, 16 bit carry lookahead low adder. 
	a4low : adder 
	generic map (
		w => 16,
		carry_logic 		=> "CLA",	-- Carry Look Ahead Logic (More Gates Used, But Less Time)
		substractor_selector	=> "NO"		-- No Just Add.
	)
	port map	(
		a => stage2p3(15 downto 0),
		b => stage2a2(15 downto 0),
		s => '0',
		ci => '0',
		result => stage2a4(15 downto 0),
		cout =>	stage2_internalCarry(1)
	);
	--! Adder 4, 16 bit carry lookahead high adder.
	a4high : adder 
	generic map (
		w => 16,
		carry_logic 		=> "CLA",	-- Carry Look Ahead Logic (More Gates Used, But Less Time)
		substractor_selector	=> "NO"		-- No Just Add.
	)
	port map	(
		a => stage2p3(31 downto 16),
		b => stage2a2(31 downto 16),
		s => '0',
		ci => stage2_internalCarry(1),
		result => stage2a4(31 downto 16),
		cout =>	open
	);	
					
	-- Incoming from opcoder.vhd signals into pipeline's stage 0.
	stage0mf00 <= m0f0;
	stage0mf01 <= m0f1;
	stage0mf10 <= m1f0;
	stage0mf11 <= m1f1;
	stage0mf20 <= m2f0;
	stage0mf21 <= m2f1;
	stage0mf30 <= m3f0;
	stage0mf31 <= m3f1;
	stage0mf40 <= m4f0;
	stage0mf41 <= m4f1;
	stage0mf50 <= m5f0;
	stage0mf51 <= m5f1;
	
	-- Signal sequencing: as the multipliers use registered output and registered input is not necessary to write the sequence of stage 0 signals to stage 1 signals.
	-- so the simplistic path is taken: simply connect stage 0 to stage 1 lines. However this would not apply for the opcode signal
	stage1p0 <= stage0p0;
	stage1p1 <= stage0p1;
	stage1p2 <= stage0p2;
	stage1p3 <= stage0p3;
	stage1p4 <= stage0p4;
	stage1p5 <= stage0p5;
	 
	
	--Outcoming to the rest of the system (by the time i wrote this i dont know where this leads to... jeje)
	cpx <= stage1a0;
	cpy <= stage1a1;
	cpz <= stage1a2;
	dp0 <= stage2a3;
	dp1 <= stage2a4;
	
	-- Looking into the design the stage 1 to stage 2 are the sequences pipe stages that must be controlled in this particular HDL.
	--! Este proceso describe la manera en que se organizan las etapas de pipe.
	--! Todas las se�ales internas en las etapas de pipe, en el momento en que la entrada rst alcanza el nivel rstMasterValue, se colocan en '0'. N�tese que, salvo stage0opcode<=stage1opcode, las se�ales que vienen desde la entrada hacia los multiplicadores en la etapa 0 y desde la salida de los multiplicadores desde la etapa0 hacia la etapa 1, no est�n siendo descritas en este proceso, la explicaci�n de es simple: Los multiplicadores que se est�n instanciado tienen registros a la entrada y la salida, permitiendo as�, registrar las entradas y registrar los productos o salidas de los  multiplicadores, hacia la etapa 1 o etapa de sumadores/restadores. 
	
	uf_seq: process (clk,rst)
	begin
		
		if rst=rstMasterValue then 
			stage0opcode	<= '0';
			stage1opcode	<= '0';
			
			stage2a2 <= (others => '0');
			stage2p3 <= (others => '0');
			stage2p2 <= (others => '0');
			stage2a0 <= (others => '0');
		
		elsif clk'event and clk = '1' then 
		
			stage2a2 <= stage1a2;
			stage2p3 <= stage1p3;
			stage2p2 <= stage1p2;
			stage2a0 <= stage1a0;
			
			-- Opcode control sequence
			stage0opcode <= opcode;
			stage1opcode <= stage0opcode;
					
		end if;
	end process uf_seq;
	
	
	
end uf_arch;
